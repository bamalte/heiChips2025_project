// SPDX-FileCopyrightText: © 2025 XXX Authors
// SPDX-License-Identifier: Apache-2.0

// Adapted from the Tiny Tapeout template

`include "alu.v"
`include "clock.v"
`include "controller.v"
`include "flags.v"
`include "ir.v"
`include "memory.v"
`include "pc.v"
`include "register.v"
`include "top.v"

`default_nettype none

module heichips25_template (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset

);

    // List all unused inputs to prevent warnings
    wire _unused = &{ena, ui_in[7:1], uio_in[7:0], uo_out/*[7:0]*/, uio_out[7:0], uio_oe[7:0]};

    top sap2_inst (
        .CLK(clk),
        .RST(~rst_n), // Active low reset
        .BUS(uio_out), // Connect only lower 8 bits of BUS to uio_out
        .A_OUT(uo_out) // Address output
    );

    
    assign uio_oe  = '1;

endmodule

